entity helloworldTB is
end entity;

-- Tip: You can input comments using "--"!

architecture sim of helloworldTB is
begin

    process is
        begin

        report "Hello World!";
        wait;

    end process;

end architecture;
